library IEEE;
use IEEE.std_logic_1164.ALL;

entity simple_vga_tb is
end simple_vga_tb;

