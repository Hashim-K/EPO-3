library IEEE;
use IEEE.std_logic_1164.ALL;

entity interr_res_tb is
end interr_res_tb;

