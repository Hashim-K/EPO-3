configuration pass_behaviour_cfg of pass is
   for behaviour
   end for;
end pass_behaviour_cfg;
