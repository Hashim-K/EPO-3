configuration clock_arch_cfg of clock is
   for arch
   end for;
end clock_arch_cfg;
