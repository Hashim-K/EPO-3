configuration eight_bit_xor_behavioural_cfg of eight_bit_xor is
   for behavioural
   end for;
end eight_bit_xor_behavioural_cfg;
