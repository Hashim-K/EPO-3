library IEEE;
use IEEE.std_logic_1164.ALL;

entity pc_high_tb is
end pc_high_tb;

