configuration eight_bit_or_behavioural_cfg of eight_bit_or is
   for behavioural
   end for;
end eight_bit_or_behavioural_cfg;
