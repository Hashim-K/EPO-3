library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of register_8bit_tb is
   component register_8bit
      port(clk     : in  std_logic;
           load    : in  std_logic;
           reset   : in  std_logic;
           data_in : in  std_logic_vector(7 downto 0);
           write   : in  std_logic;
           reg_out : out std_logic_vector(7 downto 0));
   end component;
   signal clk     : std_logic;
   signal load    : std_logic;
   signal reset   : std_logic;
   signal data_in : std_logic_vector(7 downto 0);
   signal write   : std_logic;
   signal reg_out : std_logic_vector(7 downto 0);
begin
   test: register_8bit port map (clk, load, reset, data_in, write, reg_out);
   clk <= '0' after 0 ns,
          '1' after 20 ns when clk /= '1' else '0' after 20 ns;
   load <= '0' after 0 ns,
			'1' after 40 ns,
			'0' after 80 ns,
			'1' after 120 ns,
			'0' after 200 ns;	
   reset <= '1' after 0 ns,
            '0' after 80 ns;
   data_in(0) <= '1' after 0 ns;
   data_in(1) <= '1' after 0 ns;
   data_in(2) <= '1' after 0 ns;
   data_in(3) <= '1' after 0 ns;
   data_in(4) <= '1' after 0 ns;
   data_in(5) <= '1' after 0 ns;
   data_in(6) <= '1' after 0 ns;
   data_in(7) <= '1' after 0 ns;
   write <= '0' after 0 ns,
			'1' after 80 ns,
			'0' after 120 ns,
			'1' after 160 ns;
end behaviour;

