configuration intruction_reg_synthesised_cfg of intruction_reg is
   for synthesised
   end for;
end intruction_reg_synthesised_cfg;
