configuration interr_res_behaviour_cfg of interr_res is
   for behaviour
   end for;
end interr_res_behaviour_cfg;
