library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity sprite_generator is
  port (




  -- Video output
  R : OUT std_logic;
  G : OUT std_logic;
  B : OUT std_logic
  );
end entity;

architecture arch of sprite_generator is

begin

end architecture;
