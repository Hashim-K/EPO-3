library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity instruction_register is
  port (
  clock
  );
end entity;

architecture arch of instruction_register is
begin

end architecture;
