configuration intruction_reg_tb_behaviour_sythesised_cfg of intruction_reg_tb is
   for behaviour
      for all: intruction_reg use configuration work.intruction_reg_synthesised_cfg;
      end for;
   end for;
end intruction_reg_tb_behaviour_sythesised_cfg;
