configuration eight_bit_shift_behaviour_cfg of eight_bit_shift is
   for behaviour
   end for;
end eight_bit_shift_behaviour_cfg;
