configuration interr_res_tb_behaviour_cfg of interr_res_tb is
   for behaviour
      for all: interr_res use configuration work.interr_res_behaviour_cfg;
      end for;
   end for;
end interr_res_tb_behaviour_cfg;
