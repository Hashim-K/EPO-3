library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity test is
  port (
  clock : IN std_logic;
  );
end entity;

architecture arch of test is

begin

end architecture;
