configuration intruction_reg_behaviour_cfg of intruction_reg is
   for behaviour
   end for;
end intruction_reg_behaviour_cfg;
