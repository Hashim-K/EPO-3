configuration pass_tb_behaviour_cfg of pass_tb is
   for behaviour
      for all: pass use configuration work.pass_behaviour_cfg;
      end for;
   end for;
end pass_tb_behaviour_cfg;
