configuration accumulator_tb_structural_cfg of accumulator_tb is
   for structural
      for all: accumulator use configuration work.accumulator_structural_cfg;
      end for;
   end for;
end accumulator_tb_structural_cfg;
