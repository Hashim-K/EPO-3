library ieee;

  use ieee.std_logic_1164.all;

  use ieee.numeric_std.all;


entity instruction_decoder is
  port (
      ir_in: IN STD_LOGIC_VECTOR(7 DOWNTO 0);   -- Instruction register in
      tcstate: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
      interrupt: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      ready: IN STD_LOGIC;
      r_w: OUT STD_LOGIC;
      sv: IN STD_LOGIC;
      acr : IN STD_LOGIC;
      cin : IN STD_LOGIC; -- from status register carry in
      z   : IN STD_LOGIC; -- from status register zero
      v   : IN std_logic;
      n   : IN std_logic;
      control_out: OUT STD_LOGIC_VECTOR(69 DOWNTO 0);
      s1 : IN STD_LOGIC;
      s2 : IN STD_LOGIC;
      page_crossing : OUT std_logic; -- indicate page crossing
      bcr : OUT std_logic; -- indicate branch instruction taking on
    --  ff_add: IN STD_Logic
      v1: IN STD_LOGIC
  );
end entity;

architecture arch of instruction_decoder is

-- Order of checking
  -- 1. Check CC
  -- 2. Check AAA
  -- 3. Check BBB

begin	-- TODO FIX R_W SIGNAL
	r_w <= '0';
	Control : process(tcstate, ir_in, cin) -- Fix TOM added IR, cin
	begin
case ir_in(7 downto 0) is
		when "00000000" =>
			-- Cycles:7
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000100000000000000000000000000000000110000110000001111010000000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000100000000000000000000000000000000110010110000000111000010000000000";
	--Timing: T4
elsif (tcstate(4)='0') then
--Timing: T3
	control_out<="0000110000000000000000000000000000000110010110000000111000000000000000";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0000000000000000000000000000000000000001100000000010011100101000000000";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
control_out<="0000000000000000000000000000000000000000000000000000010001100000000100";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000000000000100000010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00000001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000100001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "00000101" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000100001100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00000110" =>
			-- Cycles:5
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="1000001000000001001000000000000010000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00001000" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000110000000000000000000000000000000110000110000001111000000000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000001100000000010000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00001001" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000100001100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00001010" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000100000010000000001000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0100000100000000101000000001000000000001100000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00001101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000100001100001000000000000000000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00001110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011000000000000100";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="1000001000000001001000000000000010000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00010000" =>
			-- Cycles:4
page_crossing <= cin;
bcr <= not n;
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000001000000011100111000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0010000000000000001000000000000000000110011000000000000000000100000100";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000000000000000111100101000000000011000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "00010001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000001000000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000100001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "00010101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000011000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000100001100001000000000000000000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00010110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011000000000011000";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0010000000000000000000000000000010000000001000000000000000000000000100";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000111100100000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00011000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000100000000000000000000000000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00011001" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000001000000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000010100000000000010001000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000101000000101000000001000000100001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00011101" =>
			-- Cycles:6
page_crossing <= cin;
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
if cin = '1' then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
else
	control_out<="0000000000000000000000000010100000000000010001000000011000000000000100";
end if;
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000101000000101000000001000000100001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "00011110" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
control_out<="1000000000000000000000000000000010000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "00100000" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000100001000001100000000000000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000100000000000000000000000000000000101111000000000111000010000000000";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000100000000000000000000000000000000001110000000010111010000000000000";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000100000000000000001000000011100100000000001";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011001001100000100";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00100001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000001001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "00100100" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000001000000000011000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000100100001000000000000000000001000000001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00100101" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000001001100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00100110" =>
			-- Cycles:5
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="1000000000000000000000000000001000000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00101000" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000100001000010100000000000000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000100000000000000000000000000000000001110000000010011000000000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000100101010010010000000000000000000000000000000000000000000000001";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00101001" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000101000000101000000001000000001001100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00101010" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000100001000000000001000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0100000100000000101000000001000000000001100000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00101100" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000100100001000000000000000000001000000001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00101101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000001001100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00101110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011000000000000100";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="1000000000000000000000000000001000000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000100000000101000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00110000" =>
			-- Cycles:4
page_crossing <= cin;
bcr <= n;
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000001000000011100111000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0010000000000000001000000000000000000110011000000000000000000100000100";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000000000000000111100101000000000011000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "00110001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000001000000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000001001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "00110101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000011000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000001001100001000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00110110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011000000000011000";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0010001000000001001000000000001000000000001000000000000000000000000100";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000111100100000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00111000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000100000000000000000000000000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "00111001" =>
			-- Cycles:6
page_crossing <= cin;
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000001000000000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
if cin = '1' then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
else
	control_out<="0000000000000000000000000010100000000000010001000000011000000000000100";
end if;
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000001001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "00111101" =>
			-- Cycles:6
page_crossing <= cin;
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
if cin = '1' then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
else
	control_out<="0000000000000000000000000010100000000000010001000000011000000000000100";
end if;
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000001001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "00111110" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
control_out<="1000001000000001001000000000001000000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "01000000" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000100000000000000000000000000000000100001000010101011000000000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000100100101010010010000000000000000101111000010000011000000000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000001101000000000000001000000000100";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0000100000000000000000000000000000000100010000010000011000000000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000001100000000010000000000100000010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01000001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000010001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "01000101" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000001000000010001100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01000110" =>
			-- Cycles:5
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="1000000000000000000000000000000001000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01001000" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000100000000000000000000010000000000110000110000001111000000000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000001100000000010000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01001001" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000101000000101000000001000000010001100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01001010" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000100000001000000001000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0100000100000000101000000001000000000001100000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01001100" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000100000000000000001000000011100100000000001";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011001001100000100";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01001101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000010001101001000000000000000000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01001110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011000000000000100";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="1000000000000000000000000000000001000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000100000000101000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01010000" =>
			-- Cycles:4
page_crossing <= cin;
bcr <= not v;
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000001000000011100111000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0010000000000000001000000000000000000110011000000000000000000100000100";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000000000000000111100101000000000011000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "01010001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000001000000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000010001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "01010101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000011000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001000000000001000000010001101001000000000000000000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01010110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011000000000011000";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="1000000000000000000000000000000001000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000100000000101000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01011000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000100000000000000000000000000000000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01011001" =>
			-- Cycles:6
page_crossing <= cin;
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000001000000000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
if cin = '1' then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
else
	control_out<="0000000000000000000000000010100000000000010001000000011000000000000100";
end if;
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000101000000101000000001000000010001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "01011101" =>
			-- Cycles:6
page_crossing <= cin;
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
if cin = '1' then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
else
	control_out<="0000000000000000000000000010100000000000010001000000011000000000000100";
end if;
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000101000000101000000001000000010001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "01011110" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
control_out<="1000001000000001001000000000000001000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "01100000" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000100000000000000000000000000000000100001000010101011000000000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000001101000000000000001000000000100";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000100000000000000000000000000000000100010000010000011000000000000000";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0000000000000000000000000000000000000001100000000010000000001100000010";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000000000001000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01100001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000001000000000101100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "01100101" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000001000000000011000001000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000001000000000101100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01100110" =>
			-- Cycles:5
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="1000000000000000000000000000000100000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01101000" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000100000000000000000000100001000010100000000000000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000100000000000000000000000000000000001110000000010011000000000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="1000000000000000000000000001000000000000000000000000000000000000000001";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01101001" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000001000000000101100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01101010" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000100000100000000001000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0100000100000000101000000001000000000001100000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01101100" =>
			-- Cycles:5
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100100000000001";
--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011001001100000100";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011001001100000100";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01101101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000001000000000101100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01101110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01110000" =>
			-- Cycles:4
page_crossing <= cin;
bcr <= v;
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000001000000011100111000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0010000000000000001000000000000000000110011000000000000000000100000100";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000000000000000111100101000000000011000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "01110001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000001000000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000001000000000101100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "01110101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000011000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000001000000000101100001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01110110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011000000000011000";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="1000000000000000000000000000000100000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000100000000101000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01111000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000100000000000000000000000000000000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01111001" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000001000000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000010100000000000010001000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000001000000000101101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "01111101" =>
			-- Cycles:6
page_crossing <= cin;
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
if cin = '1' then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
else
	control_out<="0000000000000000000000000010100000000000010001000000011000000000000100";
end if;
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000001000000000101101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "01111110" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
control_out<="1000001000000001001000000000000100000000001000000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "10000001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000010000000000000000000000000111100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "10000100" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000001000000000000000000000000000000111000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10000101" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000010000000000000000000000000111000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10000110" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000010000000000000000000000000000111000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10001000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000100000000100001000000000000000100001000010000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000100000000000000001100000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10001010" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000010001000000000000000000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10001100" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000001000000000000000000010000000000111000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10001101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000010000000000000010000000000111000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10001110" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000010000000000000000010000000000111000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10010000" =>
			-- Cycles:4
page_crossing <= cin;
bcr <= not cin;
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000001000000011100111000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0010000000000000001000000000000000000110011000000000000000000100000100";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000000000000000111100101000000000011000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "10010001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000001000000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000010000000000000000000000000111100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "10010100" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000001000000000000000000010000000000111000000000011000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10010101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000010000000000000010000000000111000000000011000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10010110" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000001000000000000000100001001000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000010000000000000000010000000000111000000000011000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10011000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000001000001000000000000000000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10011001" =>
			-- Cycles:5
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000001000000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000000000000000001100000000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000010000000000000000000000000111100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "10011010" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000010000000000000000000000000010000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10011101" =>
			-- Cycles:5
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000000000000000001100000000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000010000000000000000000000000111100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "10100000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000100000000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10100001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000000001000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "10100010" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000001000000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10100100" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000100000000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10100101" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000000001000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10100110" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000001000000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10101000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000100100000000000000000000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000100000000100000000010000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10101001" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000000001000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10101010" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000001100000000000000000000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000100000000100000000010000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10101100" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000010000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000100000000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10101101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000010000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000000001000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10101110" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000010000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000001000000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10110000" =>
			-- Cycles:4
page_crossing <= cin;
bcr <= cin;
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000001000000011100111000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0010000000000000001000000000000000000110011000000000000000000100000100";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000000000000000111100101000000000011000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "10110001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000001000000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000000001000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "10110100" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000010000000000011000000000011000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000100000000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10110101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000010000000000011000000000011000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000000001000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10110110" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000001000000000000000100001001000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000010000000000011000000000011000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000001000000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10111000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0110000000000000000010000000000000000000000000000000000000000000001000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10111001" =>
			-- Cycles:6
page_crossing <= cin;
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000001000000000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
if cin = '1' then
	control_out<="0001000000000000000000000000000000000001100000000000001000000000000000";
else
	control_out<="0000000000000000000000000000000000000000010000000000011000000000000100";
end if;
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000000001000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "10111010" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000001000000000000000000000000100000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10111100" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0001000000000000000000000000000000000001100000000000001000000000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000010000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000100000000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "10111101" =>
			-- Cycles:6
page_crossing <= cin;
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
if cin = '1' then
	control_out<="0001000000000000000000000000000000000001100000000000001000000000000000";
else
	control_out<="0000000000000000000000000000000000000000010000000000011000000000000100";
end if;
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000000001000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "10111110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000001000000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0001000000000000000000000000000000000001100000000000001000000000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000010000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000100000000100000001000000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11000000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000001000000000000000000001000000000011100101000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000000000000000000000001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11000001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000100000000101000000000000000000100001000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "11000100" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000001000000000000000000001000000000011000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000100000000101000000000000000000100000000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11000101" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000001000000000011000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000100000000101000000000000000000100000000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11000110" =>
			-- Cycles:5
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="1000000100000000100000000000000000000100001000010000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000000000000000000000001000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11001000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000100000000100001000000000000000100001000001000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000100000000000000001100000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11001001" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000000000000000000000001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11001010" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000100000000100000010000000000000100001000010000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000001000000000000001100000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11001100" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000001000000000000000000011000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000000000000000100000000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11001101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000000000000000100000000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11001110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011000000000000100";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="1000001000000001000000000000000000000100001000010000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11010000" =>
			-- Cycles:4
page_crossing <= cin;
bcr <= not z;
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000001000000011100111000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0010000000000000001000000000000000000110011000000000000000000100000100";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000000000000000111100101000000000011000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "11010001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000001000000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000100000000101000000000000000000100001000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "11010101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000011000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000000000000000100000000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11010110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011000000000011000";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0000000000000000000000000000000000000010000101000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000111100100000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11011000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000010000000000000000000000000000000000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11011001" =>
			-- Cycles:6
page_crossing <= cin;
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000001000000000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
if cin = '1' then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
else
	control_out<="0000000000000000000000000010100000000000010001000000011000000000000100";
end if;
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000000000000100001101001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "11011101" =>
			-- Cycles:5
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010000000000010000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0001000000000000000000000000000000000001100000000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000100000000101000000000000000000100000000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11011110" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
control_out<="0000000000000000000000000000000000000010000101000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0100000000000000000000000000000000000001100000000000111100100000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "11100000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000000000000000000000001000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11100001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000001000000000101101000100000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "11100100" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000010000000000000000001000000000011000000000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000100000000101000000000000000000100000000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11100101" =>
			-- Cycles:3
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000001000011010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000001000000000101100000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11100110" =>
			-- Cycles:5
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="1000001000000001001000000000000000000100001000001000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="1000000000000000000000000001000000000000000000000000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11101000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000001000000001001000010000000000000100001000001000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000001000000000000001100000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11101001" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000001000000000011100101000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000101000000101000000001000000000101100000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11101010" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11101100" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000010000000000000000011000000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001000000001001000000000000000000100000000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11101101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000000010";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001001000001001000000001000000000101100000100000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11101110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000100000000000000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011000000000000100";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="1000001000000001001000000000000000000100001000001000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11110000" =>
			-- Cycles:4
page_crossing <= cin;
bcr <= z;
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000001000000011100111000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0010000000000000001000000000000000000110011000000000000000000100000100";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000000000000000111100101000000000011000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "11110001" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000001000000000000000100001001000000011100101000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011000000000011010";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001001000001001000000001000000000101101000100000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "11110101" =>
			-- Cycles:4
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000100000000000000011000000000011000000000011000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001001000001001000000001000000000101100000100000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11110110" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000000000010000000000000100001001000000000000000000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000000010000000000011000000000011000";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0000001000000001000000000000000000000010000101000000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0100000000000000000000000000000000000001100000000000111100100000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11111000" =>
			-- Cycles:2
--Timing: T0
if (tcstate(0)='0') then
control_out<="0000000000010000000000000000000000000000000000000000000000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11111001" =>
			-- Cycles:6
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000001000000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T5
	elsif (tcstate(5)='0') then
control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T0
	elsif (tcstate(0)='0') then
control_out<="0000000000000000000000000010100000000000010001000000011000000000000100";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001001000001001000000001000000100001101000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
page_crossing <= '1';
bcr <= '1';
		when "11111101" =>
			-- Cycles:6
page_crossing <= cin;
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
elsif (tcstate(3)='0') then
	control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
if cin = '1' then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
else
	control_out<="0000000000000000000000000010100000000000010001000000011000000000000100";
end if;
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000001001000001001000000001000000100001101000100000011100101000000001";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
		when "11111110" =>
			-- Cycles:7
page_crossing <= '1';
bcr <= '1';
--Timing: T2
if (tcstate(2)='0') then
	control_out<="0000000000000000000000010000000000000000001000000000011100101000000000";
--Timing: T3
	elsif (tcstate(3)='0') then
control_out<="0000000000000000001000000000000000000100000001000000011100101000000001";
	--Timing: T4
elsif (tcstate(4)='0') then
if cin = '1' then
	control_out<="0000000000000000000000000000000000000110010101000000010000000000000001";
else
	control_out<="0000000000000000000000000000000000000100010101000000010000000000000001";
end if;
--Timing: T5
	elsif (tcstate(5)='0') then
	control_out<="0001000000000000000000000010100000000001100001000000001000000000000000";
--Timing: T6
	elsif (tcstate(0)='1' and tcstate(1)='1' and tcstate(2)='1' and tcstate(3)='1' and tcstate(4)='1' and tcstate(5)='1') then
control_out<="1000001000000001000000000000000000000100001000001000000000000000000001";
--Timing: T0
	elsif (tcstate(0)='0') then
	control_out<="0100000000000000000000000000000000000001100000000000100000000000000000";
--Timing: T1
elsif (tcstate(1)='0') then
	control_out<="0000000000000000000000000000000000000000000000000000011100101000000000";
else
	control_out<="0000000000000000000000000000000000000000000000000000000000000000000000";
end if;
when OTHERS =>
control_out <= "0000000000000000000000000000000000000000000000000000000000000000000000";
end case;
end process;
end architecture;
