library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity B_input_register is
  port (
  clock
  );
end entity;

architecture arch of B_input_register is

begin

end architecture;
