library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity a_input_register is
  port (
  clock :
  );
end entity;

architecture arch of a_input_register is

begin

end architecture;
