configuration pc_low_synthesised_cfg of pc_low is
   for synthesised
   end for;
end pc_low_synthesised_cfg;
