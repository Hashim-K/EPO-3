configuration eight_bit_and_behavioural_cfg of eight_bit_and is
   for behavioural
   end for;
end eight_bit_and_behavioural_cfg;
