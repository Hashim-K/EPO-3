configuration pc_high_synthesised_cfg of pc_high is
   for synthesised
   end for;
end pc_high_synthesised_cfg;
