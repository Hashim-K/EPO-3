--Timing: T
if tcstate()='0') then
  control_out<="";
end if;
