library IEEE;
use IEEE.std_logic_1164.ALL;

entity intruction_reg_tb is
end intruction_reg_tb;

