configuration accumulator_structural_cfg of accumulator is
   for structural
      for all: register_8bit use configuration work.register_8bit_behaviour_cfg;
      end for;
   end for;
end accumulator_structural_cfg;
