library IEEE;
use IEEE.std_logic_1164.ALL;

entity pc_low_tb is

end pc_low_tb;

