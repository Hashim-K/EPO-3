configuration vga_driver_behavioural_cfg of vga_driver is
   for behavioural
   end for;
end vga_driver_behavioural_cfg;
