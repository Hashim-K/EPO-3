configuration intruction_reg_tb_behaviour_cfg of intruction_reg_tb is
   for behaviour
      for all: intruction_reg use configuration work.intruction_reg_behaviour_cfg;
      end for;
   end for;
end intruction_reg_tb_behaviour_cfg;
