configuration register_8bit_behaviour_cfg of register_8bit is
   for behaviour
   end for;
end register_8bit_behaviour_cfg;
