configuration eight_bit_adder_behaviour_cfg of eight_bit_adder is
   for behaviour
   end for;
end eight_bit_adder_behaviour_cfg;
