library IEEE;
use IEEE.std_logic_1164.ALL;

entity pass_tb is
end pass_tb;

