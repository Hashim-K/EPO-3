--Timing: T2
if (tcstate(2)='0') then
end if;
--Timing: T3
if (tcstate(3)='0') then
end if;
--Timing: T4
if (tcstate(4)='0') then
end if;
--Timing: T5
if (tcstate(5)='0') then
end if;
--Timing: T6
if (tcstate(0)='1'&tcstate(1)='1'&tcstate(2)='1'&tcstate(3)='1'&tcstate(4)='1'&tcstate(5)='1') then
end if;
--Timing: T0
if (tcstate(0)='0') then
end if;
--Timing: T1
if (tcstate(1)='0') then
end if;
