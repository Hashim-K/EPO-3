configuration a_input_register_strucutural_cfg of a_input_register is
   for strucutural
      for all: register_8bit use configuration work.register_8bit_behaviour_cfg;
      end for;
   end for;
end a_input_register_strucutural_cfg;
