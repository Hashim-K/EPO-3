configuration register_8bit_synthesised_cfg of register_8bit is
   for synthesised
   end for;
end register_8bit_synthesised_cfg;
