library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity rgb is
  port (
  clock
  );
end entity;

architecture behavioural of rgb is

begin



end architecture;
