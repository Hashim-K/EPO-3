library IEEE;
use IEEE.std_logic_1164.ALL;

entity register_8bit_tb is
end register_8bit_tb;

